library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity m4to2 is
    port(a,b,c,d: in STD_ULOGIC_VECTOR(31 downto 0);
         x, y:    out STD_ULOGIC_VECTOR(31 downto 0));
  end;
  
  architecture behav of m4to2 is
  begin
    --TODO
  end;