library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity mult is 
  port(a:   in STD_ULOGIC_VECTOR(15 downto 0);
       b:   in STD_ULOGIC_VECTOR(15 downto 0);
       y:   out STD_ULOGIC_VECTOR(31 downto 0));
end;

architecture behav of mult is 
begin
    --TODO
end;