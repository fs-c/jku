library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity CSavA is
  port(a, b, c: in STD_ULOGIC_VECTOR(31 downto 0);
       cout, s: out STD_ULOGIC_VECTOR(31 downto 0));
end;

architecture behav of CSavA is
begin
  --TODO
end; 